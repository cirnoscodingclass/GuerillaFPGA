`timescale 1ns / 1ps

module Switches_To_LEDs(
    input i_Switch_0,
    output o_LED_0
    ); 
    
    assign o_LED_0 = i_Switch_0;
endmodule
